VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

PROPERTYDEFINITIONS
  MACRO previous_effective_target_usage REAL ;
  MACRO expanded_util REAL ;
END PROPERTYDEFINITIONS

LAYER NWELL
  TYPE MASTERSLICE ;
END NWELL

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.152 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M1

LAYER VIA1
  TYPE CUT ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.152 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M2

LAYER VIA2
  TYPE CUT ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M3

LAYER VIA3
  TYPE CUT ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M4

LAYER VIA4
  TYPE CUT ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M5

LAYER VIA5
  TYPE CUT ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M6

LAYER VIA6
  TYPE CUT ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M7

LAYER VIA7
  TYPE CUT ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M8

LAYER VIA8
  TYPE CUT ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 2.432 ;
  WIDTH 0.16 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.16 WRONGDIRECTION ;" ;
END M9

LAYER VIARDL
  TYPE CUT ;
END VIARDL

LAYER MRDL
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4.864 ;
  WIDTH 2 ;
  PROPERTY LEF58_WIDTH "WIDTH 2 WRONGDIRECTION ;" ;
END MRDL

LAYER DNW
  TYPE MASTERSLICE ;
END DNW

LAYER DIFF
  TYPE MASTERSLICE ;
END DIFF

LAYER PIMP
  TYPE MASTERSLICE ;
END PIMP

LAYER NIMP
  TYPE MASTERSLICE ;
END NIMP

LAYER DIFF_18
  TYPE MASTERSLICE ;
END DIFF_18

LAYER PAD
  TYPE MASTERSLICE ;
END PAD

LAYER ESD_25
  TYPE MASTERSLICE ;
END ESD_25

LAYER SBLK
  TYPE MASTERSLICE ;
END SBLK

LAYER HVTIMP
  TYPE MASTERSLICE ;
END HVTIMP

LAYER LVTIMP
  TYPE MASTERSLICE ;
END LVTIMP

LAYER M1PIN
  TYPE MASTERSLICE ;
END M1PIN

LAYER M2PIN
  TYPE MASTERSLICE ;
END M2PIN

LAYER M3PIN
  TYPE MASTERSLICE ;
END M3PIN

LAYER M4PIN
  TYPE MASTERSLICE ;
END M4PIN

LAYER M5PIN
  TYPE MASTERSLICE ;
END M5PIN

LAYER M6PIN
  TYPE MASTERSLICE ;
END M6PIN

LAYER M7PIN
  TYPE MASTERSLICE ;
END M7PIN

LAYER M8PIN
  TYPE MASTERSLICE ;
END M8PIN

LAYER M9PIN
  TYPE MASTERSLICE ;
END M9PIN

LAYER MRDL9PIN
  TYPE MASTERSLICE ;
END MRDL9PIN

LAYER HOTNWL
  TYPE MASTERSLICE ;
END HOTNWL

LAYER DIOD
  TYPE MASTERSLICE ;
END DIOD

LAYER BJTDMY
  TYPE MASTERSLICE ;
END BJTDMY

LAYER RNW
  TYPE MASTERSLICE ;
END RNW

LAYER RMARK
  TYPE MASTERSLICE ;
END RMARK

LAYER prBoundary
  TYPE MASTERSLICE ;
END prBoundary

LAYER LOGO
  TYPE MASTERSLICE ;
END LOGO

LAYER IP
  TYPE MASTERSLICE ;
END IP

LAYER RM1
  TYPE MASTERSLICE ;
END RM1

LAYER RM2
  TYPE MASTERSLICE ;
END RM2

LAYER RM3
  TYPE MASTERSLICE ;
END RM3

LAYER RM4
  TYPE MASTERSLICE ;
END RM4

LAYER RM5
  TYPE MASTERSLICE ;
END RM5

LAYER RM6
  TYPE MASTERSLICE ;
END RM6

LAYER RM7
  TYPE MASTERSLICE ;
END RM7

LAYER RM8
  TYPE MASTERSLICE ;
END RM8

LAYER RM9
  TYPE MASTERSLICE ;
END RM9

LAYER DM1EXCL
  TYPE MASTERSLICE ;
END DM1EXCL

LAYER DM2EXCL
  TYPE MASTERSLICE ;
END DM2EXCL

LAYER DM3EXCL
  TYPE MASTERSLICE ;
END DM3EXCL

LAYER DM4EXCL
  TYPE MASTERSLICE ;
END DM4EXCL

LAYER DM5EXCL
  TYPE MASTERSLICE ;
END DM5EXCL

LAYER DM6EXCL
  TYPE MASTERSLICE ;
END DM6EXCL

LAYER DM7EXCL
  TYPE MASTERSLICE ;
END DM7EXCL

LAYER DM8EXCL
  TYPE MASTERSLICE ;
END DM8EXCL

LAYER DM9EXCL
  TYPE MASTERSLICE ;
END DM9EXCL

LAYER DIFF_25
  TYPE MASTERSLICE ;
END DIFF_25

LAYER DIFF_FM
  TYPE MASTERSLICE ;
END DIFF_FM

LAYER PO_FM
  TYPE MASTERSLICE ;
END PO_FM

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12SQ_C
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA12SQ_C

VIA VIA12BAR_C
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA12BAR_C

VIA VIA12LG_C
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG_C

VIA VIA12SQ
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA12SQ

VIA VIA12BAR
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA12BAR

VIA VIA12LG
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG

VIA VIA23SQ_C
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA23SQ_C

VIA VIA23BAR_C
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA23BAR_C

VIA VIA23LG_C
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG_C

VIA VIA23SQ
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA23SQ

VIA VIA23BAR
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA23BAR

VIA VIA23LG
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG

VIA VIA34SQ_C
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA34SQ_C

VIA VIA34BAR_C
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA34BAR_C

VIA VIA34LG_C
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG_C

VIA VIA34SQ
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA34SQ

VIA VIA34BAR
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA34BAR

VIA VIA34LG
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG

VIA VIA45SQ_C
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA45SQ_C

VIA VIA45BAR_C
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA45BAR_C

VIA VIA45LG_C
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG_C

VIA VIA45SQ
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA45SQ

VIA VIA45BAR
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA45BAR

VIA VIA45LG
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG

VIA VIA56SQ_C
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA56SQ_C

VIA VIA56BAR_C
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA56BAR_C

VIA VIA56LG_C
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG_C

VIA VIA56SQ
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA56SQ

VIA VIA56BAR
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA56BAR

VIA VIA56LG
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG

VIA VIA67SQ_C
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA67SQ_C

VIA VIA67BAR_C
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA67BAR_C

VIA VIA67LG_C
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG_C

VIA VIA67SQ
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA67SQ

VIA VIA67BAR
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA67BAR

VIA VIA67LG
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG

VIA VIA78SQ_C
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA78SQ_C

VIA VIA78BAR_C
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA78BAR_C

VIA VIA78LG_C
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG_C

VIA VIA78SQ
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA78SQ

VIA VIA78BAR
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA78BAR

VIA VIA78LG
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG

VIA VIA89_C
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.08 -0.095 0.08 0.095 ;
END VIA89_C

VIA VIA89
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.095 -0.08 0.095 0.08 ;
END VIA89

VIA VIA9RDL
  LAYER M9 ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER VIARDL ;
    RECT -1 -1 1 1 ;
  LAYER MRDL ;
    RECT -1.5 -1.5 1.5 1.5 ;
END VIA9RDL

NONDEFAULTRULE CTS_NDR_2w2s
  LAYER M2
    WIDTH 0.1 ;
    SPACING 0.1 ;
  END M2
  LAYER M3
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M3
  LAYER M4
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M4
  LAYER M5
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M5
  LAYER M6
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M6
  LAYER M7
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M7
  LAYER M8
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M8
  LAYER M9
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M9
  LAYER MRDL
    WIDTH 0.32 ;
    SPACING 0.32 ;
  END MRDL
END CTS_NDR_2w2s

NONDEFAULTRULE ndr_2w2s
  HARDSPACING ;
  LAYER M1
    WIDTH 0.1 ;
    SPACING 0.1 ;
  END M1
  LAYER M2
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M2
  LAYER M3
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M3
  LAYER M4
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M4
  LAYER M5
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M5
  LAYER M6
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M6
  LAYER M7
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M7
  LAYER M8
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M8
  LAYER M9
    WIDTH 0.32 ;
    SPACING 0.32 ;
  END M9
  LAYER MRDL
    WIDTH 4 ;
    SPACING 4 ;
  END MRDL
END ndr_2w2s

NONDEFAULTRULE ndr_2w2s_manual
  LAYER M1
    WIDTH 0.1 ;
    SPACING 0.1 ;
  END M1
  LAYER M2
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M2
  LAYER M3
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M3
  LAYER M4
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M4
  LAYER M5
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M5
  LAYER M6
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M6
  LAYER M7
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M7
  LAYER M8
    WIDTH 0.112 ;
    SPACING 0.112 ;
  END M8
  LAYER M9
    WIDTH 0.32 ;
    SPACING 0.32 ;
  END M9
  LAYER MRDL
    WIDTH 2 ;
    SPACING 2 ;
  END MRDL
END ndr_2w2s_manual

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.152 BY 1.672 ;
END unit

MACRO spi_rx
  CLASS BLOCK ;
  FOREIGN spi_rx -1.672 -1.672 ;
  ORIGIN 0 0 ;
  SIZE 23.408 BY 23.408 ;
  SYMMETRY X Y ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M5 ;
        RECT 0 8.94 0.286 8.996 ;
    END
  END clk
  PIN reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0 13.804 0.286 13.86 ;
    END
  END reset_n
  PIN sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0 10.156 0.286 10.212 ;
    END
  END sck
  PIN cs_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0 12.588 0.286 12.644 ;
    END
  END cs_n
  PIN mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0 11.372 0.286 11.428 ;
    END
  END mosi
  PIN rx_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 17.452 23.408 17.508 ;
    END
  END rx_data[7]
  PIN rx_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 16.236 23.408 16.292 ;
    END
  END rx_data[6]
  PIN rx_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 7.724 23.408 7.78 ;
    END
  END rx_data[5]
  PIN rx_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 15.02 23.408 15.076 ;
    END
  END rx_data[4]
  PIN rx_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 8.94 23.408 8.996 ;
    END
  END rx_data[3]
  PIN rx_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 13.804 23.408 13.86 ;
    END
  END rx_data[2]
  PIN rx_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 10.156 23.408 10.212 ;
    END
  END rx_data[1]
  PIN rx_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 12.588 23.408 12.644 ;
    END
  END rx_data[0]
  PIN rx_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.122 11.372 23.408 11.428 ;
    END
  END rx_valid
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
  END VSS
  OBS
    LAYER M1 SPACING 0 ;
      RECT 0 0 23.408 23.408 ;
    LAYER M2 SPACING 0 ;
      RECT 0 0 23.408 23.408 ;
    LAYER M3 SPACING 0 ;
      RECT 0 0 23.408 23.408 ;
    LAYER M4 SPACING 0 ;
      RECT 0 0 23.408 23.408 ;
    LAYER M5 SPACING 0 ;
      POLYGON 23.408 23.408 23.408 17.508 23.122 17.508 23.122 17.452 23.408 17.452 23.408 16.292 23.122 16.292 23.122 16.236 23.408 16.236 23.408 15.076 23.122 15.076 23.122 15.02 23.408 15.02 23.408 13.86 23.122 13.86 23.122 13.804 23.408 13.804 23.408 12.644 23.122 12.644 23.122 12.588 23.408 12.588 23.408 11.428 23.122 11.428 23.122 11.372 23.408 11.372 23.408 10.212 23.122 10.212 23.122 10.156 23.408 10.156 23.408 8.996 23.122 8.996 23.122 8.94 23.408 8.94 23.408 7.78 23.122 7.78 23.122 7.724 23.408 7.724 23.408 0 0 0 0 8.94 0.286 8.94 0.286 8.996 0 8.996 0 10.156 0.286 10.156 0.286 10.212 0 10.212 0 11.372 0.286 11.372 0.286 11.428 0 11.428 0 12.588 0.286 12.588 0.286 12.644 0 12.644 0 13.804 0.286 13.804 0.286 13.86 0 13.86 0 23.408 ;
    LAYER M6 SPACING 0 ;
      RECT 0 0 23.408 23.408 ;
    LAYER M7 SPACING 0 ;
      RECT 0 0 23.408 23.408 ;
    LAYER M8 SPACING 0 ;
      RECT 0 0 23.408 23.408 ;
    LAYER NWELL SPACING 0 ;
      RECT 0 0 23.408 23.408 ;
    LAYER M5 ;
      POLYGON 22.708 22.708 22.708 18.208 22.422 18.208 22.422 7.024 22.708 7.024 22.708 0.7 0.7 0.7 0.7 8.24 0.986 8.24 0.986 14.56 0.7 14.56 0.7 22.708 ;
    LAYER M1 ;
      RECT 0.6 0.6 22.808 22.808 ;
    LAYER M2 ;
      RECT 0.7 0.7 22.708 22.708 ;
    LAYER M3 ;
      POLYGON 23.007 14.47 23.007 14.41 22.897 14.41 22.897 14.412 21.1 14.412 21.1 14.468 22.897 14.468 22.897 14.47 ;
      POLYGON 0.511 13.862 0.511 13.86 2.308 13.86 2.308 13.804 0.511 13.804 0.511 13.802 0.401 13.802 0.401 13.862 ;
      POLYGON 23.007 12.342 23.007 12.282 22.897 12.282 22.897 12.284 21.1 12.284 21.1 12.34 22.897 12.34 22.897 12.342 ;
      POLYGON 0.511 8.998 0.511 8.996 2.612 8.996 2.612 8.94 0.511 8.94 0.511 8.938 0.401 8.938 0.401 8.998 ;
      RECT 0.7 0.7 22.708 22.708 ;
    LAYER M4 ;
      POLYGON 22.982 15.103 22.982 14.993 22.98 14.993 22.98 14.495 22.982 14.495 22.982 14.385 22.922 14.385 22.922 14.495 22.924 14.495 22.924 14.993 22.922 14.993 22.922 15.103 ;
      POLYGON 0.486 13.887 0.486 13.777 0.484 13.777 0.484 10.239 0.486 10.239 0.486 10.129 0.426 10.129 0.426 10.239 0.428 10.239 0.428 13.777 0.426 13.777 0.426 13.887 ;
      POLYGON 22.982 12.367 22.982 12.257 22.98 12.257 22.98 7.807 22.982 7.807 22.982 7.697 22.922 7.697 22.922 7.807 22.924 7.807 22.924 12.257 22.922 12.257 22.922 12.367 ;
      RECT 0.426 8.756 0.486 9.023 ;
      RECT 0.7 0.7 22.708 22.708 ;
    LAYER M6 ;
      RECT 0.7 0.7 22.708 22.708 ;
    LAYER M7 ;
      RECT 0.328 22.632 23.08 23.08 ;
      RECT 0.328 0.328 23.08 0.776 ;
      RECT 0.7 0.7 22.708 22.708 ;
    LAYER M8 ;
      RECT 22.632 0.328 23.08 23.08 ;
      RECT 21.016 0.328 21.24 23.08 ;
      RECT 13.72 0.328 13.944 23.08 ;
      RECT 7.64 0.328 7.864 23.08 ;
      RECT 0.328 0.328 0.776 23.08 ;
      RECT 0.7 0.7 22.708 22.708 ;
    LAYER NWELL ;
      RECT 0.23 0.23 23.178 23.178 ;
    LAYER VIA3 ;
      RECT 22.927 14.415 22.977 14.465 ;
      RECT 0.431 13.807 0.481 13.857 ;
      RECT 22.927 12.287 22.977 12.337 ;
      RECT 0.431 8.943 0.481 8.993 ;
    LAYER VIA4 ;
      RECT 22.927 15.023 22.977 15.073 ;
      RECT 0.431 10.159 0.481 10.209 ;
      RECT 0.431 8.943 0.481 8.993 ;
      RECT 22.927 7.727 22.977 7.777 ;
    LAYER VIA7 ;
      RECT 22.951 22.951 23.001 23.001 ;
      RECT 22.831 22.951 22.881 23.001 ;
      RECT 22.711 22.951 22.761 23.001 ;
      RECT 21.103 22.951 21.153 23.001 ;
      RECT 13.807 22.951 13.857 23.001 ;
      RECT 7.727 22.951 7.777 23.001 ;
      RECT 0.647 22.951 0.697 23.001 ;
      RECT 0.527 22.951 0.577 23.001 ;
      RECT 0.407 22.951 0.457 23.001 ;
      RECT 22.951 22.831 23.001 22.881 ;
      RECT 22.831 22.831 22.881 22.881 ;
      RECT 22.711 22.831 22.761 22.881 ;
      RECT 21.103 22.831 21.153 22.881 ;
      RECT 13.807 22.831 13.857 22.881 ;
      RECT 7.727 22.831 7.777 22.881 ;
      RECT 0.647 22.831 0.697 22.881 ;
      RECT 0.527 22.831 0.577 22.881 ;
      RECT 0.407 22.831 0.457 22.881 ;
      RECT 22.951 22.711 23.001 22.761 ;
      RECT 22.831 22.711 22.881 22.761 ;
      RECT 22.711 22.711 22.761 22.761 ;
      RECT 21.103 22.711 21.153 22.761 ;
      RECT 13.807 22.711 13.857 22.761 ;
      RECT 7.727 22.711 7.777 22.761 ;
      RECT 0.647 22.711 0.697 22.761 ;
      RECT 0.527 22.711 0.577 22.761 ;
      RECT 0.407 22.711 0.457 22.761 ;
      RECT 22.951 0.647 23.001 0.697 ;
      RECT 22.831 0.647 22.881 0.697 ;
      RECT 22.711 0.647 22.761 0.697 ;
      RECT 21.103 0.647 21.153 0.697 ;
      RECT 13.807 0.647 13.857 0.697 ;
      RECT 7.727 0.647 7.777 0.697 ;
      RECT 0.647 0.647 0.697 0.697 ;
      RECT 0.527 0.647 0.577 0.697 ;
      RECT 0.407 0.647 0.457 0.697 ;
      RECT 22.951 0.527 23.001 0.577 ;
      RECT 22.831 0.527 22.881 0.577 ;
      RECT 22.711 0.527 22.761 0.577 ;
      RECT 21.103 0.527 21.153 0.577 ;
      RECT 13.807 0.527 13.857 0.577 ;
      RECT 7.727 0.527 7.777 0.577 ;
      RECT 0.647 0.527 0.697 0.577 ;
      RECT 0.527 0.527 0.577 0.577 ;
      RECT 0.407 0.527 0.457 0.577 ;
      RECT 22.951 0.407 23.001 0.457 ;
      RECT 22.831 0.407 22.881 0.457 ;
      RECT 22.711 0.407 22.761 0.457 ;
      RECT 21.103 0.407 21.153 0.457 ;
      RECT 13.807 0.407 13.857 0.457 ;
      RECT 7.727 0.407 7.777 0.457 ;
      RECT 0.647 0.407 0.697 0.457 ;
      RECT 0.527 0.407 0.577 0.457 ;
      RECT 0.407 0.407 0.457 0.457 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 23.408 23.408 23.408 23.408 0 ;
  END
  PROPERTY expanded_util 0.72 ;
  PROPERTY previous_effective_target_usage 0.800000011920929 ;
END spi_rx

END LIBRARY
