VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

LAYER NWELL
  TYPE MASTERSLICE ;
END NWELL

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER CO
  TYPE CUT ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.152 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M1

LAYER VIA1
  TYPE CUT ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.152 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M2

LAYER VIA2
  TYPE CUT ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M3

LAYER VIA3
  TYPE CUT ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M4

LAYER VIA4
  TYPE CUT ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M5

LAYER VIA5
  TYPE CUT ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M6

LAYER VIA6
  TYPE CUT ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M7

LAYER VIA7
  TYPE CUT ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M8

LAYER VIA8
  TYPE CUT ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 2.432 ;
  WIDTH 0.16 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.16 WRONGDIRECTION ;" ;
END M9

LAYER VIARDL
  TYPE CUT ;
END VIARDL

LAYER MRDL
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4.864 ;
  WIDTH 2 ;
  PROPERTY LEF58_WIDTH "WIDTH 2 WRONGDIRECTION ;" ;
END MRDL

LAYER DNW
  TYPE MASTERSLICE ;
END DNW

LAYER DIFF
  TYPE MASTERSLICE ;
END DIFF

LAYER PIMP
  TYPE MASTERSLICE ;
END PIMP

LAYER NIMP
  TYPE MASTERSLICE ;
END NIMP

LAYER DIFF_18
  TYPE MASTERSLICE ;
END DIFF_18

LAYER PAD
  TYPE MASTERSLICE ;
END PAD

LAYER ESD_25
  TYPE MASTERSLICE ;
END ESD_25

LAYER SBLK
  TYPE MASTERSLICE ;
END SBLK

LAYER HVTIMP
  TYPE MASTERSLICE ;
END HVTIMP

LAYER LVTIMP
  TYPE MASTERSLICE ;
END LVTIMP

LAYER M1PIN
  TYPE MASTERSLICE ;
END M1PIN

LAYER M2PIN
  TYPE MASTERSLICE ;
END M2PIN

LAYER M3PIN
  TYPE MASTERSLICE ;
END M3PIN

LAYER M4PIN
  TYPE MASTERSLICE ;
END M4PIN

LAYER M5PIN
  TYPE MASTERSLICE ;
END M5PIN

LAYER M6PIN
  TYPE MASTERSLICE ;
END M6PIN

LAYER M7PIN
  TYPE MASTERSLICE ;
END M7PIN

LAYER M8PIN
  TYPE MASTERSLICE ;
END M8PIN

LAYER M9PIN
  TYPE MASTERSLICE ;
END M9PIN

LAYER MRDL9PIN
  TYPE MASTERSLICE ;
END MRDL9PIN

LAYER HOTNWL
  TYPE MASTERSLICE ;
END HOTNWL

LAYER DIOD
  TYPE MASTERSLICE ;
END DIOD

LAYER BJTDMY
  TYPE MASTERSLICE ;
END BJTDMY

LAYER RNW
  TYPE MASTERSLICE ;
END RNW

LAYER RMARK
  TYPE MASTERSLICE ;
END RMARK

LAYER prBoundary
  TYPE MASTERSLICE ;
END prBoundary

LAYER LOGO
  TYPE MASTERSLICE ;
END LOGO

LAYER IP
  TYPE MASTERSLICE ;
END IP

LAYER RM1
  TYPE MASTERSLICE ;
END RM1

LAYER RM2
  TYPE MASTERSLICE ;
END RM2

LAYER RM3
  TYPE MASTERSLICE ;
END RM3

LAYER RM4
  TYPE MASTERSLICE ;
END RM4

LAYER RM5
  TYPE MASTERSLICE ;
END RM5

LAYER RM6
  TYPE MASTERSLICE ;
END RM6

LAYER RM7
  TYPE MASTERSLICE ;
END RM7

LAYER RM8
  TYPE MASTERSLICE ;
END RM8

LAYER RM9
  TYPE MASTERSLICE ;
END RM9

LAYER DM1EXCL
  TYPE MASTERSLICE ;
END DM1EXCL

LAYER DM2EXCL
  TYPE MASTERSLICE ;
END DM2EXCL

LAYER DM3EXCL
  TYPE MASTERSLICE ;
END DM3EXCL

LAYER DM4EXCL
  TYPE MASTERSLICE ;
END DM4EXCL

LAYER DM5EXCL
  TYPE MASTERSLICE ;
END DM5EXCL

LAYER DM6EXCL
  TYPE MASTERSLICE ;
END DM6EXCL

LAYER DM7EXCL
  TYPE MASTERSLICE ;
END DM7EXCL

LAYER DM8EXCL
  TYPE MASTERSLICE ;
END DM8EXCL

LAYER DM9EXCL
  TYPE MASTERSLICE ;
END DM9EXCL

LAYER DIFF_25
  TYPE MASTERSLICE ;
END DIFF_25

LAYER DIFF_FM
  TYPE MASTERSLICE ;
END DIFF_FM

LAYER PO_FM
  TYPE MASTERSLICE ;
END PO_FM

VIA VIA12SQ_C
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA12SQ_C

VIA VIA12BAR_C
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA12BAR_C

VIA VIA12LG_C
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG_C

VIA VIA12SQ
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA12SQ

VIA VIA12BAR
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA12BAR

VIA VIA12LG
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG

VIA VIA23SQ_C
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA23SQ_C

VIA VIA23BAR_C
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA23BAR_C

VIA VIA23LG_C
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG_C

VIA VIA23SQ
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA23SQ

VIA VIA23BAR
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA23BAR

VIA VIA23LG
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG

VIA VIA34SQ_C
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA34SQ_C

VIA VIA34BAR_C
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA34BAR_C

VIA VIA34LG_C
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG_C

VIA VIA34SQ
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA34SQ

VIA VIA34BAR
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA34BAR

VIA VIA34LG
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG

VIA VIA45SQ_C
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA45SQ_C

VIA VIA45BAR_C
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA45BAR_C

VIA VIA45LG_C
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG_C

VIA VIA45SQ
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA45SQ

VIA VIA45BAR
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA45BAR

VIA VIA45LG
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG

VIA VIA56SQ_C
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA56SQ_C

VIA VIA56BAR_C
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA56BAR_C

VIA VIA56LG_C
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG_C

VIA VIA56SQ
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA56SQ

VIA VIA56BAR
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA56BAR

VIA VIA56LG
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG

VIA VIA67SQ_C
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA67SQ_C

VIA VIA67BAR_C
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA67BAR_C

VIA VIA67LG_C
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG_C

VIA VIA67SQ
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA67SQ

VIA VIA67BAR
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA67BAR

VIA VIA67LG
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG

VIA VIA78SQ_C
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA78SQ_C

VIA VIA78BAR_C
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA78BAR_C

VIA VIA78LG_C
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG_C

VIA VIA78SQ
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA78SQ

VIA VIA78BAR
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA78BAR

VIA VIA78LG
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG

VIA VIA89_C
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.08 -0.095 0.08 0.095 ;
END VIA89_C

VIA VIA89
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.095 -0.08 0.095 0.08 ;
END VIA89

VIA VIA9RDL
  LAYER M9 ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER VIARDL ;
    RECT -1 -1 1 1 ;
  LAYER MRDL ;
    RECT -1.5 -1.5 1.5 1.5 ;
END VIA9RDL

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.152 BY 1.672 ;
END unit

END LIBRARY
